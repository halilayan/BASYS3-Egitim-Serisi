----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Halil İbrahim Ayan
-- 
-- Create Date: 
-- Design Name: 
-- Module Name: led_animasyon - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity led_animasyon is
  Port (
        clk     : in std_logic;
        rst     : in std_logic;
        div_clk : in std_logic;
        led     : out std_logic_vector (15 downto 0)
         );
end led_animasyon;

architecture Behavioral of led_animasyon is
    type state_type is (STATE_LEFT, STATE_RIGHT);
    
    signal state            : state_type := STATE_LEFT;
    signal sequence_count   : integer range 0 to 271 := 0;
    
    type led_sequence_type is array (0 to 271) of std_logic_vector (15 downto 0);
    
    function init_led_sequence return led_sequence_type is
        variable seq : led_sequence_type;
    begin
        seq(0)   := "0000000000000001"; seq(1)   := "0000000000000010"; seq(2)   := "0000000000000100"; seq(3)   := "0000000000001000";
        seq(4)   := "0000000000010000"; seq(5)   := "0000000000100000"; seq(6)   := "0000000001000000"; seq(7)   := "0000000010000000";
        seq(8)   := "0000000100000000"; seq(9)   := "0000001000000000"; seq(10)  := "0000010000000000"; seq(11)  := "0000100000000000";
        seq(12)  := "0001000000000000"; seq(13)  := "0010000000000000"; seq(14)  := "0100000000000000"; seq(15)  := "1000000000000000";
        seq(16)  := "1000000000000001"; seq(17)  := "1000000000000010"; seq(18)  := "1000000000000100"; seq(19)  := "1000000000001000";
        seq(20)  := "1000000000010000"; seq(21)  := "1000000000100000"; seq(22)  := "1000000001000000"; seq(23)  := "1000000010000000";
        seq(24)  := "1000000100000000"; seq(25)  := "1000001000000000"; seq(26)  := "1000010000000000"; seq(27)  := "1000100000000000";
        seq(28)  := "1001000000000000"; seq(29)  := "1010000000000000"; seq(30)  := "1100000000000000"; seq(31)  := "1100000000000001"; 
        seq(32)  := "1100000000000010"; seq(33)  := "1100000000000100"; seq(34)  := "1100000000001000"; seq(35)  := "1100000000010000"; 
        seq(36)  := "1100000000100000"; seq(37)  := "1100000001000000"; seq(38)  := "1100000010000000"; seq(39)  := "1100000100000000"; 
        seq(40)  := "1100001000000000"; seq(41)  := "1100010000000000"; seq(42)  := "1100100000000000"; seq(43)  := "1101000000000000"; 
        seq(44)  := "1110000000000000"; seq(45)  := "1110000000000001"; seq(46)  := "1110000000000010"; seq(47)  := "1110000000000100"; 
        seq(48)  := "1110000000001000"; seq(49)  := "1110000000010000"; seq(50)  := "1110000000100000"; seq(51)  := "1110000001000000"; 
        seq(52)  := "1110000010000000"; seq(53)  := "1110000100000000"; seq(54)  := "1110001000000000"; seq(55)  := "1110010000000000"; 
        seq(56)  := "1110100000000000"; seq(57)  := "1111000000000000"; seq(58)  := "1111000000000001"; seq(59)  := "1111000000000010";  
        seq(60)  := "1111000000000100"; seq(61)  := "1111000000001000"; seq(62)  := "1111000000010000"; seq(63)  := "1111000000100000"; 
        seq(64)  := "1111000001000000"; seq(65)  := "1111000010000000"; seq(66)  := "1111000100000000"; seq(67)  := "1111001000000000"; 
        seq(68)  := "1111010000000000"; seq(69)  := "1111100000000000"; seq(70)  := "1111100000000001"; seq(71)  := "1111100000000010"; 
        seq(72)  := "1111100000000100"; seq(73)  := "1111100000001000"; seq(74)  := "1111100000010000"; seq(75)  := "1111100000100000"; 
        seq(76)  := "1111100001000000"; seq(77)  := "1111100010000000"; seq(78)  := "1111100100000000"; seq(79)  := "1111101000000000"; 
        seq(80)  := "1111110000000000"; seq(81)  := "1111110000000001"; seq(82)  := "1111110000000010"; seq(83)  := "1111110000000100"; 
        seq(84)  := "1111110000001000"; seq(85)  := "1111110000010000"; seq(86)  := "1111110000100000"; seq(87)  := "1111110001000000";
        seq(88)  := "1111110010000000"; seq(89)  := "1111110100000000"; seq(90)  := "1111111000000000"; seq(91)  := "1111111000000001";       
        seq(92)  := "1111111000000010"; seq(93)  := "1111111000000100"; seq(94)  := "1111111000001000"; seq(95)  := "1111111000010000";
        seq(96)  := "1111111000100000"; seq(97)  := "1111111001000000"; seq(98)  := "1111111010000000"; seq(99)  := "1111111100000000";       
        seq(100) := "1111111100000001"; seq(101) := "1111111100000010"; seq(102) := "1111111100000100"; seq(103) := "1111111100001000";
        seq(104) := "1111111100010000"; seq(105) := "1111111100100000"; seq(106) := "1111111101000000"; seq(107) := "1111111110000000";
        seq(108) := "1111111110000001"; seq(109) := "1111111110000010"; seq(110) := "1111111110000100"; seq(111) := "1111111110001000";
        seq(112) := "1111111110010000"; seq(113) := "1111111110100000"; seq(114) := "1111111111000000"; seq(115) := "1111111111000001";
        seq(116) := "1111111111000010"; seq(117) := "1111111111000100"; seq(118) := "1111111111001000"; seq(119) := "1111111111010000";
        seq(120) := "1111111111100000"; seq(121) := "1111111111100001"; seq(122) := "1111111111100010"; seq(123) := "1111111111100100";
        seq(124) := "1111111111101000"; seq(125) := "1111111111110000"; seq(126) := "1111111111110001"; seq(127) := "1111111111110010"; 
        seq(128) := "1111111111110100"; seq(129) := "1111111111111000"; seq(130) := "1111111111111001"; seq(131) := "1111111111111010";
        seq(132) := "1111111111111100"; seq(133) := "1111111111111101"; seq(134) := "1111111111111110";
        
        -- Final state: all LEDs on
        seq(135) := "1111111111111111";
        
        -- Turn-off sequence starts here
        seq(136) := "1111111111111110"; seq(137) := "1111111111111101"; seq(138) := "1111111111111100"; seq(139) := "1111111111111010";
        seq(140) := "1111111111111001"; seq(141) := "1111111111111000"; seq(142) := "1111111111110100"; seq(143) := "1111111111110010";
        seq(144) := "1111111111110001"; seq(145) := "1111111111110000"; seq(146) := "1111111111101000"; seq(147) := "1111111111100100";
        seq(148) := "1111111111100010"; seq(149) := "1111111111100001"; seq(150) := "1111111111100000"; seq(151) := "1111111111010000";
        seq(152) := "1111111111001000"; seq(153) := "1111111111000100"; seq(154) := "1111111111000010"; seq(155) := "1111111111000001";
        seq(156) := "1111111111000000"; seq(157) := "1111111110100000"; seq(158) := "1111111110010000"; seq(159) := "1111111110001000";
        seq(160) := "1111111110000100"; seq(161) := "1111111110000010"; seq(162) := "1111111110000001"; seq(163) := "1111111110000000";
        seq(164) := "1111111101000000"; seq(165) := "1111111100100000"; seq(166) := "1111111100010000"; seq(167) := "1111111100001000";
        seq(168) := "1111111100000100"; seq(169) := "1111111100000010"; seq(170) := "1111111100000001"; seq(171) := "1111111100000000";
        seq(172) := "1111111010000000"; seq(173) := "1111111001000000"; seq(174) := "1111111000100000"; seq(175) := "1111111000010000";
        seq(176) := "1111111000001000"; seq(177) := "1111111000000100"; seq(178) := "1111111000000010"; seq(179) := "1111111000000001";
        seq(180) := "1111111000000000"; seq(181) := "1111110100000000"; seq(182) := "1111110010000000"; seq(183) := "1111110001000000";
        seq(184) := "1111110000100000"; seq(185) := "1111110000010000"; seq(186) := "1111110000001000"; seq(187) := "1111110000000100";
        seq(188) := "1111110000000010"; seq(189) := "1111110000000001"; seq(190) := "1111110000000000"; seq(191) := "1111101000000000";
        seq(192) := "1111100100000000"; seq(193) := "1111100010000000"; seq(194) := "1111100001000000"; seq(195) := "1111100000100000";
        seq(196) := "1111100000010000"; seq(197) := "1111100000001000"; seq(198) := "1111100000000100"; seq(199) := "1111100000000010";
        seq(200) := "1111100000000001"; seq(201) := "1111100000000000"; seq(202) := "1111010000000000"; seq(203) := "1111001000000000";
        seq(204) := "1111000100000000"; seq(205) := "1111000010000000"; seq(206) := "1111000001000000"; seq(207) := "1111000000100000";
        seq(208) := "1111000000010000"; seq(209) := "1111000000001000"; seq(210) := "1111000000000100"; seq(211) := "1111000000000010";
        seq(212) := "1111000000000001"; seq(213) := "1111000000000000"; seq(214) := "1110100000000000"; seq(215) := "1110010000000000";
        seq(216) := "1110001000000000"; seq(217) := "1110000100000000"; seq(218) := "1110000010000000"; seq(219) := "1110000001000000";
        seq(220) := "1110000000100000"; seq(221) := "1110000000010000"; seq(222) := "1110000000001000"; seq(223) := "1110000000000100";
        seq(224) := "1110000000000010"; seq(225) := "1110000000000001"; seq(226) := "1110000000000000"; seq(227) := "1101000000000000";
        seq(228) := "1100100000000000"; seq(229) := "1100010000000000"; seq(230) := "1100001000000000"; seq(231) := "1100000100000000";
        seq(232) := "1100000010000000"; seq(233) := "1100000001000000"; seq(234) := "1100000000100000"; seq(235) := "1100000000010000";
        seq(236) := "1100000000001000"; seq(237) := "1100000000000100"; seq(238) := "1100000000000010"; seq(239) := "1100000000000001";
        seq(240) := "1100000000000000"; seq(241) := "1010000000000000"; seq(242) := "1001000000000000"; seq(243) := "1000100000000000";
        seq(244) := "1000010000000000"; seq(245) := "1000001000000000"; seq(246) := "1000000100000000"; seq(247) := "1000000010000000";
        seq(248) := "1000000001000000"; seq(249) := "1000000000100000"; seq(250) := "1000000000010000"; seq(251) := "1000000000001000";
        seq(252) := "1000000000000100"; seq(253) := "1000000000000010"; seq(254) := "1000000000000001"; seq(255) := "1000000000000000";
        seq(256) := "0100000000000000"; seq(257) := "0010000000000000"; seq(258) := "0001000000000000"; seq(259) := "0000100000000000";
        seq(260) := "0000010000000000"; seq(261) := "0000001000000000"; seq(262) := "0000000100000000"; seq(263) := "0000000010000000";
        seq(264) := "0000000001000000"; seq(265) := "0000000000100000"; seq(266) := "0000000000010000"; seq(267) := "0000000000001000";
        seq(268) := "0000000000000100"; seq(269) := "0000000000000010"; seq(270) := "0000000000000001"; seq(271) := "0000000000000000";
        return seq;
    end function;
    
    signal led_sequence : led_sequence_type := init_led_sequence;

begin

    process(clk)
        begin
            if rising_edge(clk) then
                if rst = '1' then
                    sequence_count <= 0;
                    state <= STATE_LEFT;
                elsif div_clk = '1' then
                    case state is
                        when STATE_LEFT =>
                            if sequence_count < 135 then
                                sequence_count <= sequence_count + 1;
                            else 
                                state <= STATE_RIGHT;
                            end if;
                        
                        when STATE_RIGHT =>
                            if sequence_count < 271 then 
                                sequence_count <= sequence_count +1;
                            else
                                state <= STATE_LEFT;
                                sequence_count <= 0;
                            end if;
                    end case; 
                
                end if;
            
            end if;
    end process;
    
    led <= led_sequence(sequence_count);


end Behavioral;
